--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.VECTOR_STANDARD.ALL;

--A package containing declarations of constant parameter sets
--Of Elliptic Curve Domain Parameters.
package ECC_STANDARD is

----------------------------------------------------
-----------Declare types of generic size!-----------
----------------------------------------------------

type ECC_Parameters_521 is array (0 to 5) of STD_LOGIC_VECTOR(520 downto 0);
type ECC_Parameters_384 is array (0 to 5) of STD_LOGIC_VECTOR(383 downto 0);
type ECC_Parameters_256 is array (0 to 5) of STD_LOGIC_VECTOR(255 downto 0);
type ECC_Parameters_224 is array (0 to 5) of STD_LOGIC_VECTOR(223 downto 0);
type ECC_Parameters_192 is array (0 to 5) of STD_LOGIC_VECTOR(191 downto 0);
type ECC_Parameters_160 is array (0 to 5) of STD_LOGIC_VECTOR(159 downto 0);
type ECC_Parameters_128 is array (0 to 5) of STD_LOGIC_VECTOR(127 downto 0);
type ECC_Parameters_112 is array (0 to 5) of STD_LOGIC_VECTOR(111 downto 0);
type ECC_Parameters_5 is array (0 to 5) of STD_LOGIC_VECTOR(4 downto 0);

----------------------------------
-----------Naming model-----------
----------------------------------

----Curve_Name
--constant Curve_Name : ECC_Parameters_BitLength := (
--X"Hex String", --Prime
--X"Hex String", --A
--X"Hex String", --B
--X"Hex String", --GX
--X"Hex String", --GY
--X"Hex String");--N

-------------------------------------
-----------List of Curves!-----------
-------------------------------------

--SECp521r1
constant SECp521r1 : ECC_Parameters_521 := (
"1" & X"FF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF", --Prime
"1" & X"FF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFC", --A
"0" & X"51_953E_B961_8E1C_9A1F_929A_21A0_B685_40EE_A2DA_725B_99B3_15F3_B8B4_8991_8EF1_09E1_5619_3951_EC7E_937B_1652_C0BD_3BB1_BF07_3573_DF88_3D2C_34F1_EF45_1FD4_6B50_3F00", --B
"0" & X"C6_858E_06B7_0404_E9CD_9E3E_CB66_2395_B442_9C64_8139_053F_B521_F828_AF60_6B4D_3DBA_A14B_5E77_EFE7_5928_FE1D_C127_A2FF_A8DE_3348_B3C1_856A_429B_F97E_7E31_C2E5_BD66", --GX
"1" & X"18_3929_6A78_9A3B_C004_5C8A_5FB4_2C7D_1BD9_98F5_4449_579B_4468_17AF_BD17_273E_662C_97EE_7299_5EF4_2640_C550_B901_3FAD_0761_353C_7086_A272_C240_88BE_9476_9FD1_6650", --GY
"1" & X"FF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFA_5186_8783_BF2F_966B_7FCC_0148_F709_A5D0_3BB5_C9B8_899C_47AE_BB6F_B71E_9138_6409");--N

--SECp384r1
constant SECp384r1 : ECC_Parameters_384 := (
X"FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFE_FFFF_FFFF_0000_0000_0000_0000_FFFF_FFFF", --Prime
X"FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFE_FFFF_FFFF_0000_0000_0000_0000_FFFF_FFFC", --A
X"B331_2FA7_E23E_E7E4_988E_056B_E3F8_2D19_181D_9C6E_FE81_4112_0314_088F_5013_875A_C656_398D_8A2E_D19D_2A85_C8ED_D3EC_2AEF", --B
X"AA87_CA22_BE8B_0537_8EB1_C71E_F320_AD74_6E1D_3B62_8BA7_9B98_59F7_41E0_8254_2A38_5502_F25D_BF55_296C_3A54_5E38_7276_0AB7", --GX
X"3617_DE4A_9626_2C6F_5D9E_98BF_9292_DC29_F8F4_1DBD_289A_147C_E9DA_3113_B5F0_B8C0_0A60_B1CE_1D7E_819D_7A43_1D7C_90EA_0E5F", --GY
X"FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_C763_4D81_F437_2DDF_581A_0DB2_48B0_A77A_ECEC_196A_CCC5_2973");--N

--SECp256r1
constant SECp256r1 : ECC_Parameters_256 := (
X"FFFF_FFFF_0000_0001_0000_0000_0000_0000_0000_0000_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF", --Prime
X"FFFF_FFFF_0000_0001_0000_0000_0000_0000_0000_0000_FFFF_FFFF_FFFF_FFFF_FFFF_FFFC", --A
X"5AC6_35D8_AA3A_93E7_B3EB_BD55_7698_86BC_651D_06B0_CC53_B0F6_3BCE_3C3E_27D2_604B", --B
X"6B17_D1F2_E12C_4247_F8BC_E6E5_63A4_40F2_7703_7D81_2DEB_33A0_F4A1_3945_D898_C296", --GX
X"4FE3_42E2_FE1A_7F9B_8EE7_EB4A_7C0F_9E16_2BCE_3357_6B31_5ECE_CBB6_4068_37BF_51F5", --GY
X"FFFF_FFFF_0000_0000_FFFF_FFFF_FFFF_FFFF_BCE6_FAAD_A717_9E84_F3B9_CAC2_FC63_2551");--N

--SECp256k1
constant SECp256k1 : ECC_Parameters_256 := (
X"FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFE_FFFF_FC2F", --Prime
X"0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000", --A
X"0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0007", --B
X"79BE_667E_F9DC_BBAC_55A0_6295_CE87_0B07_029B_FCDB_2DCE_28D9_59F2_815B_16F8_1798", --GX
X"483A_DA77_26A3_C465_5DA4_FBFC_0E11_08A8_FD17_B448_A685_5419_9C47_D08F_FB10_D4B8", --GY
X"FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFE_BAAE_DCE6_AF48_A03B_BFD2_5E8C_D036_4141");--N

--SECp224k1: Not implemented, N is longer in bitlength than the prime.

--SECp224r1
constant SECp224r1 : ECC_Parameters_224 := (
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_00000000_00000000_00000001", --Prime
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFE_FFFFFFFF_FFFFFFFF_FFFFFFFE", --A
X"B4050A85_0C04B3AB_F5413256_5044B0B7_D7BFD8BA_270B3943_2355FFB4", --B
X"B70E0CBD_6BB4BF7F_321390B9_4A03C1D3_56C21122_343280D6_115C1D21", --GX
X"BD376388_B5F723FB_4C22DFE6_CD4375A0_5A074764_44D58199_85007E34", --GY
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFF16A2_E0B8F03E_13DD2945_5C5C2A3D");--N

--SECp192k1
constant SECp192k1 : ECC_Parameters_192 := (
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFE_FFFFEE37", --Prime
X"00000000_00000000_00000000_00000000_00000000_00000000", --A
X"00000000_00000000_00000000_00000000_00000000_00000003", --B
X"DB4FF10E_C057E9AE_26B07D02_80B7F434_1DA5D1B1_EAE06C7D", --GX
X"9B2F2F6D_9C5628A7_844163D0_15BE8634_4082AA88_D95E2F9D", --GY
X"FFFFFFFF_FFFFFFFF_FFFFFFFE_26F2FC17_0F69466A_74DEFD8D");--N

--SECp192r1
constant SECp192r1 : ECC_Parameters_192 := (
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFE_FFFFFFFF_FFFFFFFF", --Prime
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFE_FFFFFFFF_FFFFFFFC", --A
X"64210519_E59C80E7_0FA7E9AB_72243049_FEB8DEEC_C146B9B1", --B
X"188DA80E_B03090F6_7CBF20EB_43A18800_F4FF0AFD_82FF1012", --GX
X"07192B95_FFC8DA78_631011ED_6B24CDD5_73F977A1_1E794811", --GY
X"FFFFFFFF_FFFFFFFF_FFFFFFFF_99DEF836_146BC9B1_B4D22831");--N

----SECp160k1: Not implemented, N is longer in bitlength than the prime.
----SECp160r1: Not implemented, N is longer in bitlength than the prime.
----SECp160r2: Not implemented, N is longer in bitlength than the prime.

--SECp128r1
constant SECp128r1 : ECC_Parameters_128 := (
X"FFFFFFFD_FFFFFFFF_FFFFFFFF_FFFFFFFF", --Prime
X"FFFFFFFD_FFFFFFFF_FFFFFFFF_FFFFFFFC", --A
X"E87579C1_1079F43D_D824993C_2CEE5ED3", --B
X"161FF752_8B899B2D_0C28607C_A52C5B86", --GX
X"CF5AC839_5BAFEB13_C02DA292_DDED7A83", --GY
X"FFFFFFFE_00000000_75A30D1B_9038A115");--N

--SECp128r2
constant SECp128r2 : ECC_Parameters_128 := (
X"FFFFFFFD_FFFFFFFF_FFFFFFFF_FFFFFFFF", --Prime
X"D6031998_D1B3BBFE_BF59CC9B_BFF9AEE1", --A
X"5EEEFCA3_80D02919_DC2C6558_BB6D8A5D", --B
X"7B6AA5D8_5E572983_E6FB32A7_CDEBC140", --GX
X"27B6916A_894D3AEE_7106FE80_5FC34B44", --GY
X"3FFFFFFF_7FFFFFFF_BE002472_0613B5A3");--N

--SECp112r1
constant SECp112r1 : ECC_Parameters_112 := (
X"DB7C_2ABF_62E3_5E66_8076_BEAD_208B", --Prime
X"DB7C_2ABF_62E3_5E66_8076_BEAD_2088", --A
X"659E_F8BA_0439_16EE_DE89_1170_2B22", --B
X"0948_7239_995A_5EE7_6B55_F9C2_F098", --GX
X"A89C_E5AF_8724_C0A2_3E0E_0FF7_7500", --GY
X"DB7C_2ABF_62E3_5E76_28DF_AC65_61C5");--N

--SECp112r2
constant SECp112r2 : ECC_Parameters_112 := (
X"DB7C_2ABF_62E3_5E66_8076_BEAD_208B", --Prime
X"6127_C24C_05F3_8A0A_AAF6_5C0E_F02C", --A
X"51DE_F181_5DB5_ED74_FCC3_4C85_D709", --B
X"4BA3_0AB5_E892_B4E1_649D_D092_8643", --GX
X"ADCD_46F5_882E_3747_DEF3_6E95_6E97", --GY
X"36DF_0AAF_D8B8_D759_7CA1_0520_D04B");--N

--M17
constant M17 : ECC_Parameters_5 := (
"10001", --Prime
"00010", --A
"00010", --B
"00111", --GX
"00110", --GY
"10011");--N

-----------------------------------------------------------------------------
-----------Legacy Curves, left here for use by older library files-----------
-----------------------------------------------------------------------------

--SECp256r1 (non-typed)
constant Prime_NISTsecp256r1 : STD_LOGIC_VECTOR (255 downto 0) := X"FFFF_FFFF_0000_0001_0000_0000_0000_0000_0000_0000_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF";
constant Prime_NISTsecp256r1_2Compliment : STD_LOGIC_VECTOR (255 downto 0) := X"0000_0000_FFFF_FFFE_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_0000_0000_0000_0000_0000_0001";
constant A_NISTsecp256r1 : STD_LOGIC_VECTOR (255 downto 0) := X"FFFF_FFFF_0000_0001_0000_0000_0000_0000_0000_0000_FFFF_FFFF_FFFF_FFFF_FFFF_FFFC";
constant B_NISTsecp256r1 : STD_LOGIC_VECTOR (255 downto 0) := X"5AC6_35D8_AA3A_93E7_B3EB_BD55_7698_86BC_651D_06B0_CC53_B0F6_3BCE_3C3E_27D2_604B";
constant GX_NISTsecp256r1 : STD_LOGIC_VECTOR (255 downto 0) := X"6B17_D1F2_E12C_4247_F8BC_E6E5_63A4_40F2_7703_7D81_2DEB_33A0_F4A1_3945_D898_C296";
constant GY_NISTsecp256r1 : STD_LOGIC_VECTOR (255 downto 0) := X"4FE3_42E2_FE1A_7F9B_8EE7_EB4A_7C0F_9E16_2BCE_3357_6B31_5ECE_CBB6_4068_37BF_51F5";
constant N_NISTsecp256r1 : STD_LOGIC_VECTOR (255 downto 0) := X"FFFFFFFF_00000000_FFFFFFFF_FFFFFFFF_BCE6FAAD_A7179E84_F3B9CAC2_FC632551";
--M17 (non-typed)
constant Prime_M17 : STD_LOGIC_VECTOR (4 downto 0) := "10001";
constant Prime_M17_2Compliment : STD_LOGIC_VECTOR (4 downto 0) := "01111";
constant A_M17 : STD_LOGIC_VECTOR (4 downto 0) := "00010";
constant B_M17 : STD_LOGIC_VECTOR (4 downto 0) := "00010";
constant GX_M17 : STD_LOGIC_VECTOR (4 downto 0) := "00111";
constant GY_M17 : STD_LOGIC_VECTOR (4 downto 0) := "00110";

end ECC_STANDARD;

package body ECC_STANDARD is
 
end ECC_STANDARD;
